.circuit
V1 n1 GND dc 7
V2 n1 n2 dc 5
V3 n2 GND dc 2  #loops of voltage sources
.end
