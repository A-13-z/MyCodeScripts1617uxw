.circuit
V1 1 GND dc 5
V2 1 2 dc 9
R1 2 GND 1
V3 1 3 dc 7
R2 3 GND 2
.end