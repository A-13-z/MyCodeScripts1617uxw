.circuit
I1 GND n1 3
.end

#single current source